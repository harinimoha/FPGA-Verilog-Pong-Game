module Motion_Ball (
    input clock,
    input reset,
    input start_game,
    input [15:0] paddle1_Y,
    input [15:0] paddle2_Y,
    output reg [15:0] Ball_X,
    output reg [15:0] Ball_Y,
    output reg [15:0] Vx,
    output reg [15:0] Vy
);

    // Parameters for screen resolution, ball size, and initial velocities
    parameter SCREEN_WIDTH = 640;
    parameter SCREEN_HEIGHT = 480;
    parameter BALL_SIZE = 10;
    parameter INITIAL_VX = 0;
    parameter INITIAL_VY = 0;

    // These are the states in which the ball directions could be in (six possible directions)
    localparam UP = 3'b000;
    localparam DOWN = 3'b001;
    localparam LEFT_UP = 3'b010;
    localparam LEFT_DOWN = 3'b011;
    localparam RIGHT_UP = 3'b100;
    localparam RIGHT_DOWN = 3'b101;

    // These would temporarily hold updated values for use by the game to ensure that the motion of the ball is continuous. 
    reg [2:0] direction;
    reg [15:0] next_Ball_X;
    reg [15:0] next_Ball_Y;
    reg [15:0] next_Vx;
    reg [15:0] next_Vy;

    always @(posedge clock or posedge reset) 
    begin
        if (reset) 
            begin
            // Initialize ball position and velocities
            Ball_X <= SCREEN_WIDTH / 2 - BALL_SIZE / 2;
            Ball_Y <= SCREEN_HEIGHT / 2 - BALL_SIZE / 2;

            Vx <= INITIAL_VX;
            Vy <= INITIAL_VY;

            direction <= UP;
            end
 
            else if (start_game) 
            begin
            // Updating ball position based on current velocities
            next_Ball_X = Ball_X + Vx;
            next_Ball_Y = Ball_Y + Vy;

            // Checking for collision with paddles and updating velocities

            case (direction)
                UP: 
					 begin

                    // Check if the ball collided with the top wall
                    if (next_Ball_Y <= 0) 
                        begin
                        direction <= DOWN; // Collide with upper wall and move downwards
                        end

                    // Check if the ball collided with paddle 1
                    else if ((next_Ball_X <= 20) && (next_Ball_Y >= paddle1_Y) && (next_Ball_Y < paddle1_Y + 80)) 
			           begin
                        direction <= RIGHT_DOWN;        // Move diagonally downward towards Paddle 2
                    end

                    // Check if the ball collided with paddle 2
                    else if ((next_Ball_X >= SCREEN_WIDTH - 20 - BALL_SIZE) && (next_Ball_Y >= paddle2_Y) && (next_Ball_Y < paddle2_Y + 80)) 
			           begin
                        direction <= LEFT_DOWN;        // Move diagonally downward towards Paddle 1
                    end

                 end

                DOWN: 
		    begin
                    // Check if the ball collided with the bottom wall and move upward if it does. 
                    if (next_Ball_Y >= SCREEN_HEIGHT - BALL_SIZE) 
                        begin
                        direction <= UP; // Reflect upward
                        end

                    // Check if the ball collided with paddle 1 
                    else if ((next_Ball_X <= 20) && (next_Ball_Y >= paddle1_Y) && (next_Ball_Y < paddle1_Y + 80)) 
			begin
                        direction <= RIGHT_UP; // Move diagonally upward towards Paddle 2
                        end

                    // Check if the ball collided with paddle 2
                    else if ((next_Ball_X >= SCREEN_WIDTH - 20 - BALL_SIZE) && (next_Ball_Y >= paddle2_Y) && (next_Ball_Y < paddle2_Y + 80))
		        begin
                        direction <= LEFT_UP; // Move diagonally upward towards Paddle 1
                        end
                    end

                LEFT_UP: 
                    begin

                    // Check if the ball collided with Paddle 1
                    if ((next_Ball_X <= 20) && (next_Ball_Y >= paddle1_Y) && (next_Ball_Y < paddle1_Y + 80)) 
                    	begin
                        direction <= RIGHT_UP; // Reflect upward
                    	end

                    // Check if the ball  collided with Paddle 2
                    else if ((next_Ball_X >= SCREEN_WIDTH - 20 - BALL_SIZE) && (next_Ball_Y >= paddle2_Y) && (next_Ball_Y < paddle2_Y + 80)) 
                    	begin
                        direction <= LEFT_UP; // Reflect upward
                    	end

                    // Check if the ball collided with the top wall
                    else if (next_Ball_Y <= 0) 
			begin
                        direction <= LEFT_DOWN; // Move diagonally downward towards Paddle 1
                    	end

                    end

                LEFT_DOWN: 
	            begin
                    // Check if the ball coincided with Paddle 1
                    if ((next_Ball_X <= 20) && (next_Ball_Y >= paddle1_Y) && (next_Ball_Y < paddle1_Y + 80)) begin
                        direction <= RIGHT_DOWN;       // Reflect downward
                    end

                    // Check if paddle coincided with Paddle 2
                    else if ((next_Ball_X >= SCREEN_WIDTH - 20 - BALL_SIZE) && (next_Ball_Y >= paddle2_Y) && (next_Ball_Y < paddle2_Y + 80)) begin
                        direction <= LEFT_DOWN;        // Reflect downward
                    end

                    // Check if paddle coincided with bottom wall
                    else if (next_Ball_Y >= SCREEN_HEIGHT - BALL_SIZE) 
						  begin
                        direction <= LEFT_UP;          // Move diagonally upward towards Paddle 1
                    end

                end

                RIGHT_UP: 
                    begin
                    // Check if the ball collided with Paddle 1
                    if ((next_Ball_X <= 20) && (next_Ball_Y >= paddle1_Y) && (next_Ball_Y < paddle1_Y + 80)) begin
                        direction <= RIGHT_UP; // Reflect upward
                    end

                    // Check if the ball collided with Paddle 2
                    else if ((next_Ball_X >= SCREEN_WIDTH - 20 - BALL_SIZE) && (next_Ball_Y >= paddle2_Y) && (next_Ball_Y < paddle2_Y + 80)) begin
                        direction <= LEFT_UP; // Reflect upward
                    end

                    // Check if the ball collided with top wall
                    else if (next_Ball_Y <= 0) begin
                        direction <= RIGHT_DOWN; // Move diagonally downward towards Paddle 2
                    end
                end
                RIGHT_DOWN: begin
                    // Check for collision with Paddle 1
                    if ((next_Ball_X <= 20) && (next_Ball_Y >= paddle1_Y) && (next_Ball_Y < paddle1_Y + 80)) 
		    begin
                        direction <= RIGHT_DOWN; // Reflect downward
                    end

                    // Check for collision with Paddle 2
                    else if ((next_Ball_X >= SCREEN_WIDTH - 20 - BALL_SIZE) && (next_Ball_Y >= paddle2_Y) && (next_Ball_Y < paddle2_Y + 80)) 
                    begin
                        direction <= LEFT_DOWN; // Reflect downward
                    end

                    // Check for collision with bottom wall
                    else if (next_Ball_Y >= SCREEN_HEIGHT - BALL_SIZE) 
		    begin
                        direction <= RIGHT_UP; // Move diagonally upward towards Paddle 2
                    end
                end

                default: 
                    begin
                    	Ball_X <= SCREEN_WIDTH / 2 - BALL_SIZE / 2;
            		Ball_Y <= SCREEN_HEIGHT / 2 - BALL_SIZE / 2;
                    end
            endcase

            // Updated velocities based on new locations 
            case (direction)
                UP: 
                begin
                    next_Vx = 0;
                    next_Vy = -2;
                end

                DOWN: 
                begin
                    next_Vx = 0;
                    next_Vy = 2;
                end

                LEFT_UP: 
                begin
                    next_Vx = -2;
                    next_Vy = -2;
                end

                LEFT_DOWN: 
                begin
                    next_Vx = -2;
                    next_Vy = 2;
                end

                RIGHT_UP: 
                begin
                    next_Vx = 1;
                    next_Vy = -1;
                end

                RIGHT_DOWN: 
		begin
                    next_Vx = 1;
                    next_Vy = 1;
                end

                default: 
                begin
		    next_Vx = 0;
                    next_Vy = 0;   
                end

            endcase

        end

        // Now, the state variable will be updated accordingly as the game runs. 

        Ball_X <= next_Ball_X;
        Ball_Y <= next_Ball_Y;
        Vx <= next_Vx;
        Vy <= next_Vy;

    end

endmodule